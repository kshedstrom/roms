netcdf clm_ts {

dimensions:
	xi_rho = 130 ;
	xi_u = 129 ;
	xi_v = 130 ;
	eta_rho = 130 ;
	eta_u = 130 ;
	eta_v = 129 ;
	s_rho = 20 ;
	s_w = 21 ;
	tracer = 2 ;
	temp_time = 12 ;
	salt_time = 12 ;

variables:
        char spherical ;
                spherical:long_name = "grid type logical switch" ;
                spherical:flag_values = "T, F" ;
                spherical:flag_meanings = "spherical Cartesian" ;
        int Vtransform ;
                Vtransform:long_name = "vertical terrain-following transformation equation" ;
        int Vstretching ;
                Vstretching:long_name = "vertical terrain-following stretching function" ;
        double theta_s ;
                theta_s:long_name = "S-coordinate surface control parameter" ;
                theta_s:units = "nondimensional" ;
        double theta_b ;
                theta_b:long_name = "S-coordinate bottom control parameter" ;
                theta_b:units = "nondimensional" ;
        double Tcline ;
                Tcline:long_name = "S-coordinate surface/bottom layer width" ;
                Tcline:units = "meter" ;
        double hc ;
                hc:long_name = "S-coordinate parameter, critical depth" ;
                hc:units = "meter" ;
        double s_rho(s_rho) ;
                s_rho:long_name = "S-coordinate at RHO-points" ;
                s_rho:valid_min = -1. ;
                s_rho:valid_max = 0. ;
                s_rho:positive = "up" ;
                s_rho:standard_name = "ocean_s_coordinate_g1" ;
                s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
        double s_w(s_w) ;
                s_w:long_name = "S-coordinate at W-points" ;
                s_w:valid_min = -1. ;
                s_w:valid_max = 0. ;
                s_w:positive = "up" ;
                s_w:standard_name = "ocean_s_coordinate_g1" ;
                s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
        double Cs_r(s_rho) ;
                Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
                Cs_r:valid_min = -1. ;
                Cs_r:valid_max = 0. ;
        double Cs_w(s_w) ;
                Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
                Cs_w:valid_min = -1. ;
                Cs_w:valid_max = 0. ;
        double h(eta_rho, xi_rho) ;
                h:long_name = "bathymetry at RHO-points" ;
                h:units = "meter" ;
                h:coordinates = "lon_rho lat_rho" ;
        double lon_rho(eta_rho, xi_rho) ;
                lon_rho:long_name = "longitude of RHO-points" ;
                lon_rho:units = "degree_east" ;
                lon_rho:standard_name = "longitude" ;
        double lat_rho(eta_rho, xi_rho) ;
                lat_rho:long_name = "latitude of RHO-points" ;
                lat_rho:units = "degree_north" ;
                lat_rho:standard_name = "latitude" ;
	double temp_time(temp_time) ;
		temp_time:long_name = "time for potential temperature" ;
		temp_time:units = "day" ;
		temp_time:cycle_length = 360. ;
	double salt_time(salt_time) ;
		salt_time:long_name = "time for salinity" ;
		salt_time:units = "day" ;
		salt_time:cycle_length = 360. ;
	float temp(temp_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "temp_time" ;
                temp:coordinates = "lon_rho lat_rho s_rho temp_time" ;
	float salt(salt_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "salt_time" ;
                salt:coordinates = "lon_rho lat_rho s_rho salt_time" ;

// global attributes:
		:type = "CLIMATOLOGY file" ;
		:title = "Levitus One-Degree Monthly T-S Climatology (1994) - DAMEE #4" ;
		:out_file = "damee4_Lclm.nc" ;
		:grd_file = "damee4_grid_a.nc" ;
		:history = "Version 4.0  , Tuesday - March 21, 2000 - 4:47:16 PM" ;

}
