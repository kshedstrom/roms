netcdf s4dvar_std_f {

dimensions:
        xi_rho = 62 ;
        xi_u = 61 ;
        xi_v = 62 ;
        xi_psi = 61 ;
        eta_rho = 62 ;
        eta_u = 62 ;
        eta_v = 61 ;
        eta_psi = 61 ;
        N = 30 ;
        s_rho = 30 ;
        s_w = 30 ;
        ocean_time = UNLIMITED ; // (0 currently)

variables:
        char spherical ;
                spherical:long_name = "grid type logical switch" ;
                spherical:flag_values = "T, F" ;
                spherical:flag_meanings = "spherical Cartesian" ;
        int Vtransform ;
                Vtransform:long_name = "vertical terrain-following transformation equation" ;
        int Vstretching ;
                Vstretching:long_name = "vertical terrain-following stretching function" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
		theta_s:units = "nondimensional" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
		theta_b:units = "nondimensional" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
                s_rho:positive = "up" ;
                s_rho:standard_name = "ocean_s_coordinate_g1" ;
                s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
                s_w:positive = "up" ;
                s_w:standard_name = "ocean_s_coordinate_g1" ;
                s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
        double h(eta_rho, xi_rho) ;
                h:long_name = "bathymetry at RHO-points" ;
                h:units = "meter" ;
                h:coordinates = "lon_rho lat_rho" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
                lon_rho:standard_name = "longitude" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
                lat_rho:standard_name = "latitude" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
                lon_u:standard_name = "longitude" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
                lat_u:standard_name = "latitude" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
                lon_v:standard_name = "longitude" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
                lat_v:standard_name = "latitude" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "averaged time since initialization" ;
		ocean_time:units = "seconds since 2006-01-01 00:00:00" ;
		ocean_time:calendar = "365.25_day" ;
        double sustr(ocean_time, eta_u, xi_u) ;
                sustr:long_name = "surface u-momentum stress standard deviation" ;
                sustr:units = "newton meter-2" ;
                sustr:time = "ocean_time" ;
                sustr:coordinates = "lat_u lon_u ocean_time" ;
        double svstr(ocean_time, eta_v, xi_v) ;
                svstr:long_name = "surface v-momentum stress standard deviation" ;
                svstr:units = "newton meter-2" ;
                svstr:time = "ocean_time" ;
                svstr:coordinates = "lat_v lon_v ocean_time" ;
        double shflux(ocean_time, eta_rho, xi_rho) ;
                shflux:long_name = "surface net heat flux standard deviation" ;
                shflux:units = "watt meter-2" ;
                shflux:negative_value = "upward flux, cooling" ;
                shflux:positive_value = "downward flux, heating" ;
                shflux:time = "ocean_time" ;
                shflux:coordinates = "lat_rho lon_rho ocean_time" ;
        double swflux(ocean_time, eta_rho, xi_rho) ;
                swflux:long_name = "surface net freshwater flux (E-P) standard deviation" ;
                swflux:units = "meter second-1" ;
                swflux:negative_value = "upward flux, freshening (net precipitation)" ;
                swflux:positive_value = "downward flux, salting (net evaporation)" ;
                swflux:time = "ocean_time" ;
                swflux:coordinates = "lat_rho lon_rho ocean_time" ;

// global attributes:
		:type = "ROMS/TOMS 4DVAR surface forcing error covariance standard deviation" ;
		:Conventions = "CF-1.0" ;
		:title = "ROMS/TOMS 3.0 - Shallow Water 2006 Experiment, Coarse Grid" ;
}
