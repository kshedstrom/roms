netcdf s4dvar_std_f {

dimensions:
        xi_rho = 62 ;
        xi_u = 61 ;
        xi_v = 62 ;
        xi_psi = 61 ;
        eta_rho = 62 ;
        eta_u = 62 ;
        eta_v = 61 ;
        eta_psi = 61 ;
        N = 30 ;
        s_rho = 30 ;
        s_w = 30 ;
        ocean_time = UNLIMITED ; // (0 currently)

variables:
	char spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:option_T = "spherical" ;
		spherical:option_F = "Cartesian" ;
        double theta_s ;
                theta_s:long_name = "S-coordinate surface control parameter" ;
        double theta_b ;
                theta_b:long_name = "S-coordinate bottom control parameter" ;
        double Tcline ;
                Tcline:long_name = "S-coordinate surface/bottom layer width" ;
                Tcline:units = "meter" ;
        double hc ;
                hc:long_name = "S-coordinate parameter, critical depth" ;
                hc:units = "meter" ;
        double s_rho(s_rho) ;
                s_rho:long_name = "S-coordinate at RHO-points" ;
                s_rho:valid_min = -1. ;
                s_rho:valid_max = 0. ;
                s_rho:standard_name = "ocean_s_coordinate" ;
                s_rho:formula_terms = "s: s_rho eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
                s_rho:field = "s_rho, scalar" ;
        double s_w(s_w) ;
                s_w:long_name = "S-coordinate at W-points" ;
                s_w:valid_min = -1. ;
                s_w:valid_max = 0. ;
                s_w:standard_name = "ocean_s_coordinate" ;
                s_w:formula_terms = "s: s_w eta: zeta depth: h a: theta_s b: theta_b depth_c: hc" ;
                s_w:field = "s_w, scalar" ;
        double Cs_r(s_rho) ;
                Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
                Cs_r:valid_min = -1. ;
                Cs_r:valid_max = 0. ;
                Cs_r:field = "Cs_r, scalar" ;
        double Cs_w(s_w) ;
                Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
                Cs_w:valid_min = -1. ;
                Cs_w:valid_max = 0. ;
                Cs_w:field = "Cs_w, scalar" ;
        double h(eta_rho, xi_rho) ;
                h:long_name = "bathymetry at RHO-points" ;
                h:units = "meter" ;
                h:coordinates = "lon_rho lat_rho" ;
                h:field = "bath, scalar" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:field = "lon_rho, scalar" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:field = "lat_rho, scalar" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
		lon_u:field = "lon_u, scalar" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
		lat_u:field = "lat_u, scalar" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
		lon_v:field = "lon_v, scalar" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
		lat_v:field = "lat_v, scalar" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between XI-axis and EAST" ;
		angle:units = "radians" ;
		angle:coordinates = "lat_rho lon_rho" ;
		angle:field = "angle, scalar" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:option_0 = "land" ;
		mask_rho:option_1 = "water" ;
		mask_rho:coordinates = "lat_rho lon_rho" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:option_0 = "land" ;
		mask_u:option_1 = "water" ;
		mask_u:coordinates = "lat_u lon_u" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:option_0 = "land" ;
		mask_v:option_1 = "water" ;
		mask_v:coordinates = "lat_v lon_v" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "averaged time since initialization" ;
		ocean_time:units = "seconds since 2006-01-01 00:00:00" ;
		ocean_time:calendar = "365.25_day" ;
		ocean_time:field = "time, scalar, series" ;
        double sustr(ocean_time, eta_u, xi_u) ;
                sustr:long_name = "surface u-momentum stress standard deviation" ;
                sustr:units = "newton meter-2" ;
                sustr:time = "ocean_time" ;
                sustr:coordinates = "lat_u lon_u ocean_time" ;
                sustr:field = "surface u-momentum stress, scalar, series" ;
        double svstr(ocean_time, eta_v, xi_v) ;
                svstr:long_name = "surface v-momentum stress standard deviation" ;
                svstr:units = "newton meter-2" ;
                svstr:time = "ocean_time" ;
                svstr:coordinates = "lat_v lon_v ocean_time" ;
                svstr:field = "surface v-momentum stress, scalar, series" ;
        double shflux(ocean_time, eta_rho, xi_rho) ;
                shflux:long_name = "surface net heat flux standard deviation" ;
                shflux:units = "watt meter-2" ;
                shflux:negative_value = "upward flux, cooling" ;
                shflux:positive_value = "downward flux, heating" ;
                shflux:time = "ocean_time" ;
                shflux:coordinates = "lat_rho lon_rho ocean_time" ;
                shflux:field = "surface heat flux, scalar, series" ;
        double swflux(ocean_time, eta_rho, xi_rho) ;
                swflux:long_name = "surface net freshwater flux (E-P) standard deviation" ;
                swflux:units = "meter second-1" ;
                swflux:negative_value = "upward flux, freshening (net precipitation)" ;
                swflux:positive_value = "downward flux, salting (net evaporation)" ;
                swflux:time = "ocean_time" ;
                swflux:coordinates = "lat_rho lon_rho ocean_time" ;
                swflux:field = "surface net freshwater flux, scalar, series" ;
// global attributes:
		:type = "ROMS/TOMS 4DVAR surface forcing error covariance standard deviation file" ;
		:Conventions = "CF-1.0" ;
		:title = "ROMS/TOMS 3.0 - Shallow Water 2006 Experiment, Coarse Grid" ;
}
